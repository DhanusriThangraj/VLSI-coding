// 1. 1 22 333 4444 55555 4444 333 22 1 display this sequence in diamond shape 
// design code
module diamond_shape;
    initial begin
  $display("1      ");
  $display("22      ");
  $display("333      ");
  $display("4444      ");
  $display("55555      ");
  $display("4444      ");
  $display("333      ");
  $display("22      ");
  $display("1      ");
    end
endmodule

// output
1      
22      
333      
4444      
55555      
4444      
333      
22      
1 
