// design code
module carry_look_ahead_carry_generator(
  input wire [3:0]a,
  input wire [3:0]b,
  input wire cin,

  output reg cout
   );
  wire [3:0] G;
  wire [3:0] P;
  wire [3:1] c;
  
  assign G=a&b;
  assign P=a^b;
  
  assign c[1]=G[0]|(P[0]&cin);
  assign c[2]=G[1]|(P[1]&G[0])|(P[1]&P[0]&cin);
  assign c[3]=G[2]|(P[2]&G[1])|(P[2]&P[1]&G[0])|(P[2]&P[1]&P[0]&cin);
  assign cout=G[3]|(P[3]&G[2])|(P[3]&P[2]&G[1])|(P[3]&P[2]&P[1]&G[0])|(P[3]&P[2]&P[1]&P[0]&cin);
  
endmodule

// testbench
module carry_look_ahead_carry_generator_tb;
  reg [3:0]a;
  reg [3:0]b;
  reg cin;
  
  wire cout;
   
  carry_look_ahead_carry_generator uut (a,b,cin,cout);
  
  initial begin
    $display ("Time\ta\tb\tcin\tcout\t");
    $monitor("%0t\t%b\t%b\t%b\t%b",$time,a,b,cin,cout);
    
    #1; a=4'b0010; b=4'b0101; cin=1;
    #5; a=4'b1010; b=4'b0101; cin=0;
    #5; a=4'b1110; b=4'b0111; cin=1;
    #5; a=4'b0011; b=4'b1101; cin=0;
    #5; a=4'b1010; b=4'b0111; cin=1;
    #2; $finish;
  end 
endmodule
