module top_module(
    input clk,
    input areset,    // Asynchronous reset to OFF
    input j,
    input k,
    output out); //  

    parameter OFF=0, ON=1; 
    reg state, next_state;

    always @(*) begin
        case(state)
        ON:begin next_state=k?OFF:ON; end      
        OFF:begin next_state=j?ON:OFF; end
       endcase
    end

    always @(posedge clk, posedge areset) begin
        if (areset) 
            state<=OFF;
        else
            state<= next_state;
    end
    assign out = (state == ON)?1'b1:1'b0;
endmodule
